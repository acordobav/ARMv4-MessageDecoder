module romtb();


endmodule 